library ieee;
use ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;
entity instrMemory is
 port ( 
   Addr : in  std_logic_vector(3 downto 0);
   C    : out std_logic_vector(31 downto 0));
end instrMemory;

architecture arch1 of instrMemory is
signal rom_addr: std_logic_vector(3 downto 0);
  
  -- add $4, $5, $6 = 6
  type instr_array is array (0 to 15) of std_logic_vector (31 downto 0);
  constant instrmem: instr_array := ( 
	"11111111111111111111111111111111",
	"00000000000000000000000000000000",
	"11111111111111111111111111111111",
	"00000000000000000000000000000000",
	"11111111111111111111111111111111",
	"00000000101001100010000000100000",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111",
	"11111111111111111111111111111111");
begin
  C <= instrmem(to_integer(unsigned(Addr)));
end arch1;

